module ascii_pixel(
    char,
    xpos,
    ypos,
    white
    );

    input [6:0] char;
    input [1:0] xpos;
    input [2:0] ypos;

    output white;

    wire [2:0] pixels [127:0] [5:0];

    assign pixel = pixels[char][ypos][xpos];

const unsigned char ASCII[256][6] = 
{{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},/*A*/{0b01000000,0b10100000,0b11100000,0b10100000,0b10100000,0b00000000},/*B*/{0b11000000,0b10100000,0b11000000,0b10100000,0b11000000,0b00000000},/*C*/{0b01100000,0b10000000,0b10000000,0b10000000,0b01100000,0b00000000},/*D*/{0b11000000,0b10100000,0b10100000,0b10100000,0b11000000,0b00000000},/*E*/{0b11100000,0b10000000,0b11000000,0b10000000,0b11100000,0b00000000},/*F*/{0b11100000,0b10000000,0b11000000,0b10000000,0b10000000,0b00000000},/*G*/{0b01100000,0b10000000,0b10100000,0b10100000,0b01100000,0b00000000},/*H*/{0b10100000,0b10100000,0b11100000,0b10100000,0b10100000,0b00000000},/*I*/{0b11100000,0b01000000,0b01000000,0b01000000,0b11100000,0b00000000},/*J*/{0b00100000,0b00100000,0b00100000,0b10100000,0b01000000,0b00000000},/*K*/{0b10100000,0b10100000,0b11000000,0b10100000,0b10100000,0b00000000},/*L*/{0b10000000,0b10000000,0b10000000,0b10000000,0b11100000,0b00000000},/*M*/{0b10100000,0b11100000,0b10100000,0b10100000,0b10100000,0b00000000},/*N*/{0b11000000,0b10100000,0b10100000,0b10100000,0b10100000,0b00000000},/*O*/{0b11100000,0b10100000,0b10100000,0b10100000,0b11100000,0b00000000},/*P*/{0b11000000,0b10100000,0b11000000,0b10000000,0b10000000,0b00000000},/*Q*/{0b01000000,0b10100000,0b10100000,0b11100000,0b01100000,0b00000000},/*R*/{0b11000000,0b10100000,0b11000000,0b10100000,0b10100000,0b00000000},/*S*/{0b01100000,0b10000000,0b01000000,0b00100000,0b11000000,0b00000000},/*T*/{0b11100000,0b01000000,0b01000000,0b01000000,0b01000000,0b00000000},/*U*/{0b10100000,0b10100000,0b10100000,0b10100000,0b11100000,0b00000000},/*V*/{0b10100000,0b10100000,0b10100000,0b01000000,0b01000000,0b00000000},/*W*/{0b10100000,0b10100000,0b10100000,0b11100000,0b10100000,0b00000000},/*X*/{0b10100000,0b10100000,0b01000000,0b10100000,0b10100000,0b00000000},/*Y*/{0b10100000,0b10100000,0b01000000,0b01000000,0b01000000,0b00000000},/*Z*/{0b11100000,0b00100000,0b01000000,0b10000000,0b11100000,0b00000000},/* 
*/{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},/* 
*/{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},/* 
*/{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},/* 
*/{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},/* 
*/{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},/* 
*/{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},/*a*/{0b00000000,0b01100000,0b10100000,0b10100000,0b01100000,0b00000000},/*b*/{0b10000000,0b11000000,0b10100000,0b10100000,0b11000000,0b00000000},/*c*/{0b00000000,0b01100000,0b10000000,0b10000000,0b01100000,0b00000000},/*d*/{0b00100000,0b01100000,0b10100000,0b10100000,0b01100000,0b00000000},/*e*/{0b00000000,0b01000000,0b10100000,0b11000000,0b01100000,0b00000000},/*f*/{0b01100000,0b10000000,0b11000000,0b10000000,0b10000000,0b00000000},/*g*/{0b00000000,0b01100000,0b10100000,0b01100000,0b00100000,0b11000000},/*h*/{0b10000000,0b11000000,0b10100000,0b10100000,0b10100000,0b00000000},/*i*/{0b01000000,0b00000000,0b01000000,0b01000000,0b01000000,0b00000000},/*j*/{0b00100000,0b00000000,0b00100000,0b00100000,0b10100000,0b01000000},/*k*/{0b10000000,0b10000000,0b10100000,0b11000000,0b10100000,0b00000000},/*l*/{0b11000000,0b01000000,0b01000000,0b01000000,0b01000000,0b00000000},/*m*/{0b00000000,0b10100000,0b11100000,0b10100000,0b10100000,0b00000000},/*n*/{0b00000000,0b11000000,0b10100000,0b10100000,0b10100000,0b00000000},/*o*/{0b00000000,0b01000000,0b10100000,0b10100000,0b01000000,0b00000000},/*p*/{0b00000000,0b11000000,0b10100000,0b10100000,0b11000000,0b10000000},/*q*/{0b00000000,0b01100000,0b10100000,0b10100000,0b01100000,0b00100000},/*r*/{0b00000000,0b10100000,0b11000000,0b10000000,0b10000000,0b00000000},/*s*/{0b00000000,0b01100000,0b11000000,0b00100000,0b11000000,0b00000000},/*t*/{0b10000000,0b11100000,0b10000000,0b10000000,0b01100000,0b00000000},/*u*/{0b00000000,0b10100000,0b10100000,0b10100000,0b01100000,0b00000000},/*v*/{0b00000000,0b10100000,0b10100000,0b10100000,0b01000000,0b00000000},/*w*/{0b00000000,0b10100000,0b10100000,0b11100000,0b10100000,0b00000000},/*x*/{0b00000000,0b10100000,0b01000000,0b01000000,0b10100000,0b00000000},/*y*/{0b00000000,0b10100000,0b10100000,0b10100000,0b01000000,0b10000000},/*z*/{0b00000000,0b11100000,0b01000000,0b10000000,0b11100000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000},{0b00000000,0b00000000,0b00000000,0b00000000,0b00000000,0b00000000}};
endmodule
